module BCD(temp, Display);
	input [3:0] temp;
	output [0:6] Display;
	
	assign Display [0:6] = (temp[3:0] == 4'b0000) ? 7'b0000001: //0
							(temp[3:0] == 4'b0001) ? 7'b1001111: //1
							(temp[3:0] == 4'b0010) ? 7'b0010010: //2
							(temp[3:0] == 4'b0011) ? 7'b0000110: //3
							(temp[3:0] == 4'b0100) ? 7'b1001100: //4
							(temp[3:0] == 4'b0101) ? 7'b0100100: //5
							(temp[3:0] == 4'b0110) ? 7'b0100000: //6
							(temp[3:0] == 4'b0111) ? 7'b0001111: //7
							(temp[3:0] == 4'b1000) ? 7'b0000000: 7'b0000100; //8 else 9
endmodule